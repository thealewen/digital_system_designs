module toplevel(
	input logic [9:0] switches,
	input logic Clk, Run, Continue,
	output logic [9:0] LED,
	output logic [6:0] HEX0, HEX1, HEX2, HEX3
);



endmodule
