//8-bit serial logic processor

module Processor_8 (input logic	Clk,		// Clock signal for processor
											Flag,		// Extend functions of the 2 buttons on FPGA
											Reset_Execute,		// Reset (Flag = 0) signal to initialize controller to start
																	// Execute (Flag = 1) start processor execution
											LoadA_LoadB,			// Loads Register A (Flag = 0) or B (Flag = 1)
							input logic	[7:0] Din,		//data
							input logic [2:0] F,			// function select
							input logic [1:0] R,			// router select
							output logic [3:0]  LED,     // DEBUG
							output logic [7:0]  Aval,    // DEBUG
													Bval,    // DEBUG
							output logic [6:0]  AhexL,
													AhexU,
													BhexL,
													BhexU			);
													
	 logic Res_Ex_SH, LDA_LDB_SH
	 logic [2:0] F_S;
	 logic [1:0] R_S;
	 logic Ld_A, Ld_B, newA, newB, outputA, outputB, bitA, bitB, Shift_En,
	       F_A_B;
	 logic [7:0] A, B, Din_S;
	 
	 
	 //We can use the "assign" statement to do simple combinational logic
	 assign Aval = A;
	 assign Bval = B;
	 assign LED = {Execute_SH,LoadA_SH,LoadB_SH,Reset_SH}; //Concatenate is a common operation in HDL
	 
	 //Instantiation of modules here
	 register_unit_8    reg_unit_8 (
                        .Clk(Clk),
                        .Reset(Reset_SH),
                        .Ld_A, //note these are inferred assignments, because of the existence a logic variable of the same name
                        .Ld_B,
                        .Shift_En,
                        .D(Din_S),
                        .A_In(newA),
                        .B_In(newB),
                        .A_out(outputA),
                        .B_out(outputB),
                        .A(A),
                        .B(B) );
		router           router (
								.R(R_S),
                        .A_In(bitA),
                        .B_In(bitB),
                        .A_Out(newA),
                        .B_Out(newB),
                        .F_A_B );
		compute_8         compute_unit_8 (
								.F(F_S),
                        .A_In(outputA),
                        .B_In(outputB),
                        .A_Out(bitA),
                        .B_Out(bitB),
                        .F_A_B );
		control          control_unit (
                        .Clk(Clk),
                        .Reset(Reset_SH),
                        .LoadA(LoadA_SH),
                        .LoadB(LoadB_SH),
                        .Execute(Execute_SH),
                        .Shift_En,
                        .Ld_A,
                        .Ld_B );
		HexDriver        HexAL (
                        .In0(A[3:0]),
                        .Out0(AhexL) );
	 HexDriver        HexBL (
                        .In0(B[3:0]),
                        .Out0(BhexL) );
								
	 HexDriver        HexAU (
                        .In0(A[7:4]),
                        .Out0(AhexU) );	
	 HexDriver        HexBU (
                       .In0(B[7:4]),
                        .Out0(BhexU) );
								

	sync button_sync[3:0] (Clk, {~Reset, ~LoadA, ~LoadB, ~Execute}, {Reset_SH, LoadA_SH, LoadB_SH, Execute_SH});
	  sync Din_sync[3:0] (Clk, Din, Din_S);
	  sync F_sync[2:0] (Clk, F, F_S);
	  sync R_sync[1:0] (Clk, R, R_S);
	 
endmodule
		